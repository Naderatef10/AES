/* key expansion module used to generate the required key each round for the add round key operation in the AES operation
the key expansion mainly depends on the round number which is generated from the counter module, 
the enable_key_expansion is generated from the top level controller to enable key expansion each round
key expansion is bypassed in the initial round as the input key is used so the module will act as a buffer between input and output
*/

module key_expansion (
input wire clk,
input wire rst, 
input wire [3:0] round_number, /*input from the counter module*/
input wire bypass, /*input from top level controller to bypass the input in the initial round*/
input wire enable_key_expansion, /*input from top level controller to enable the operations every round*/

/*input old keys from the previous round*/
input wire [7:0] K0,
input wire [7:0] K1,
input wire [7:0] K2,
input wire [7:0] K3,
input wire [7:0] K4,
input wire [7:0] K5,
input wire [7:0] K6,
input wire [7:0] K7,
input wire [7:0] K8,
input wire [7:0] K9,
input wire [7:0] K10,
input wire [7:0] K11,
input wire [7:0] K12,
input wire [7:0] K13,
input wire [7:0] K14,
input wire [7:0] K15,


/*new 16 bytes keys after performing the expansion process*/
output reg [7:0] K0_new,
output reg [7:0] K1_new,
output reg [7:0] K2_new,
output reg [7:0] K3_new,
output reg [7:0] K4_new,
output reg [7:0] K5_new,
output reg [7:0] K6_new,
output reg [7:0] K7_new,
output reg [7:0] K8_new,
output reg [7:0] K9_new,
output reg [7:0] K10_new,
output reg [7:0] K11_new,
output reg [7:0] K12_new,
output reg [7:0] K13_new,
output reg [7:0] K14_new,
output reg [7:0] K15_new
);

/******************************intermediate signals used in the module*****************/
reg [15:0] R_conn; /*Signal needed in key expansion and it's value change according to the round number it will be implemented as a LUT*/

/*substituted bytes as the last column in the key matrix will be shifted and then subsituted using sbox matrix from the fips standard*/
wire [7:0] K_13_sub;
wire [7:0] K_14_sub;
wire [7:0] K_15_sub;
wire [7:0] K_12_sub;



/*combinational logic output to separate the combinational logic from the sequential logic*/
reg [7:0] K0_new_comb;
reg [7:0] K1_new_comb;
reg [7:0] K2_new_comb;
reg [7:0] K3_new_comb;
reg [7:0] K4_new_comb;
reg [7:0] K5_new_comb;
reg [7:0] K6_new_comb;
reg [7:0] K7_new_comb;
reg [7:0] K8_new_comb;
reg [7:0] K9_new_comb;
reg [7:0] K10_new_comb;
reg [7:0] K11_new_comb;
reg [7:0] K12_new_comb;
reg [7:0] K13_new_comb;
reg [7:0] K14_new_comb;
reg [7:0] K15_new_comb;






/*substiuting the last column of the key matrix which will be used to calculate the new first column of the key matrix*/
sbox s1(K13,K_13_sub);
sbox s2(K14,K_14_sub);
sbox s3(K15,K_15_sub);
sbox s4(K12,K_12_sub);

/*generate R_conn signal according to the round number, the values are extracted from the fips standard*/
always @(*) begin
    
    case (round_number)

        4'd1: R_conn = 16'h01;

        4'd2: R_conn = 16'h02;

        4'd3: R_conn = 16'h04;

        4'd4: R_conn = 16'h08;

        4'd5: R_conn = 16'h10;

        4'd6: R_conn = 16'h20;

        4'd7: R_conn = 16'h40;

        4'd8: R_conn = 16'h80;

        4'd9: R_conn = 16'h1B;

        4'd10: R_conn = 16'h36;
        default : R_conn = 0;
        
    endcase
end
/*combinational logic*/
always @(*) begin
    /*if bypass is enabled the output will be the same as the input*/
    if(bypass)begin
            K0_new_comb= K0;
            K1_new_comb= K1;
            K2_new_comb= K2;
            K3_new_comb= K3;
            K4_new_comb= K4;
            K5_new_comb=K5;
            K6_new_comb=K6;
            K7_new_comb=K7;
            K8_new_comb=K8;
            K9_new_comb=K9;
            K10_new_comb=K10;
            K11_new_comb=K11;
            K12_new_comb=K12;
            K13_new_comb=K13;
            K14_new_comb=K14;
            K15_new_comb=K15;                 
    end
    /*if the key expansion is enabled (once each round)*/
    else if (enable_key_expansion) begin
        /*  k0 k4 k8 k12
            k1 k5 k9 k13
            k2 k6 k10 k14
            k3 k7 k11 k15
        */

        /*first column of the key matrix*/  
            K0_new_comb = (K0 ^ K_13_sub ^ R_conn);    /*first byte is generated from xoring the old byte with the substituted byte and rconn
            after performing one cyclic shift*/
            /*  k13 -> K13_sub (output of sbox)
                k14 -> k14_sub (output of sbox)
                k15 -> k15_sub (output of sbox)
                k12 -> k12_sub (output of sbox)
            */
            /*xoring between the old byte and the corresponding byte after shifting and substituting*/
            K1_new_comb =  (K1^K_14_sub);
            K2_new_comb = (K2^K_15_sub);
            K3_new_comb = (K3^K_12_sub);

            /*second column of the key matrix*/
            /*generated by xoring the previous (from previous round) second column with the new first column (current round) of the key matrix*/
            K4_new_comb = K4 ^ K0_new_comb;
            K5_new_comb = K5 ^ K1_new_comb;
            K6_new_comb = K6 ^ K2_new_comb;
            K7_new_comb = K7 ^ K3_new_comb;
            /*third column of the key matrix*/
            /*generated by xoring the previous (from previous round) third column with the new second column (current round) of the key matrix*/
            K8_new_comb = K8 ^ K4_new_comb;
            K9_new_comb = K9 ^ K5_new_comb;
            K10_new_comb = K10 ^K6_new_comb;
            K11_new_comb = K11 ^ K7_new_comb;
            /*fourth column of the key matrix*/
            /*generated by xoring the previous (from previous round) fourth column with the new third column (current round) of the key matrix*/
            K12_new_comb = K12 ^ K8_new_comb;
            K13_new_comb = K13 ^ K9_new_comb;
            K14_new_comb = K14 ^ K10_new_comb;
            K15_new_comb = K15 ^ K11_new_comb;

        
    end
    else begin /*if not bypassed or enabled bypass*/
            K0_new_comb= K0;
            K1_new_comb= K1;
            K2_new_comb= K2;
            K3_new_comb= K3;
            K4_new_comb= K4;
            K5_new_comb=K5;
            K6_new_comb=K6;
            K7_new_comb=K7;
            K8_new_comb=K8;
            K9_new_comb=K9;
            K10_new_comb=K10;
            K11_new_comb=K11;
            K12_new_comb=K12;
            K13_new_comb=K13;
            K14_new_comb=K14;
            K15_new_comb=K15;
    end


end
/*registering the combinational logic*/

always @(posedge clk , negedge rst) begin

        if(!rst)begin
            K0_new<=0;
            K1_new<=0;
            K2_new<=0;
            K3_new<=0;
            K4_new<=0;
            K5_new<=0;
            K6_new<=0;
            K7_new<=0;
            K8_new<=0;
            K9_new<=0;
            K10_new<=0;
            K11_new<=0;
            K12_new<=0;
            K13_new<=0;
            K14_new<=0;
            K15_new<=0;
        end
        else begin
            K0_new<=K0_new_comb;
            K1_new<=K1_new_comb;
            K2_new<=K2_new_comb;
            K3_new<=K3_new_comb;
            K4_new<=K4_new_comb;
            K5_new<=K5_new_comb;
            K6_new<=K6_new_comb;
            K7_new<=K7_new_comb;
            K8_new<=K8_new_comb;
            K9_new<=K9_new_comb;
            K10_new<=K10_new_comb;
            K11_new<=K11_new_comb;
            K12_new<=K12_new_comb;
            K13_new<=K13_new_comb;
            K14_new<=K14_new_comb;
            K15_new<=K15_new_comb;

        end
end

    
endmodule